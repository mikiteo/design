--core top, will be later